/*priya branch check*/
`include "../ALU/ALU.v"
`include "../data_memory/data_memory.v"
`include "../Registers/Register.v"
module top(input clk,reset);

reg PC
