module control(input )